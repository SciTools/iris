dimensions:
	projection_y_coordinate = UNLIMITED ; // (3 currently)
	projection_x_coordinate = 4 ;
variables:
	int64 air_pressure_anomaly(projection_y_coordinate, projection_x_coordinate) ;
		air_pressure_anomaly:standard_name = "air_pressure_anomaly" ;
		air_pressure_anomaly:grid_mapping = "transverse_mercator" ;
	int transverse_mercator ;
		transverse_mercator:grid_mapping_name = "transverse_mercator" ;
		transverse_mercator:longitude_of_central_meridian = -2. ;
		transverse_mercator:latitude_of_projection_origin = 49. ;
		transverse_mercator:false_easting = -400000. ;
		transverse_mercator:false_northing = 100000. ;
		transverse_mercator:scale_factor_at_central_meridian = 0.9996012717 ;
	int64 projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	int64 projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
}
