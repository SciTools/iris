dimensions:
	depth = 20 ;
	time = 16 ;
variables:
	float m__s44i101(depth, time) ;
		m__s44i101:_FillValue = 9.96921e+36f ;
		m__s44i101:um_stash_source = "m??s44i101" ;
		m__s44i101:cell_methods = "time: mean (interval: 24 hour)" ;
	float depth(depth) ;
		depth:axis = "Z" ;
		depth:units = "m" ;
		depth:standard_name = "depth" ;
		depth:positive = "down" ;
	float time(time) ;
		time:axis = "T" ;
		time:units = "days since 0000-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;

// global attributes:
		:source = "Data from Met Office Unified Model" ;
		:Conventions = "CF-1.5" ;
}
