dimensions:
	bnds = 2 ;
	latitude = 94 ;
	longitude = 128 ;
variables:
	float sea_surface_height_above_geoid(latitude, longitude) ;
		sea_surface_height_above_geoid:_FillValue = -1.e+30f ;
		sea_surface_height_above_geoid:standard_name = "sea_surface_height_above_geoid" ;
		sea_surface_height_above_geoid:units = "m" ;
		sea_surface_height_above_geoid:grid_mapping = "latitude_longitude" ;
		sea_surface_height_above_geoid:coordinates = "forecast_period forecast_reference_time time" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	double forecast_period ;
		forecast_period:bounds = "forecast_period_bnds" ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	double forecast_period_bnds(bnds) ;
	double forecast_reference_time ;
		forecast_reference_time:units = "hours since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "360_day" ;
	double time ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(bnds) ;

// global attributes:
		:Conventions = "CF-1.5" ;
}
