dimensions:
	Mesh2_edge_N_faces = 2 ;
	Mesh2_edge_N_nodes = 2 ;
	Mesh2_face_N_edges = 4 ;
	Mesh2_face_N_faces = 4 ;
	Mesh2_face_N_nodes = 4 ;
	Mesh2_layers = 10 ;
	nMesh2_edge = 7 ;
	nMesh2_face = 2 ;
	nMesh2_node = 6 ;
variables:
	int Mesh2 ;
		Mesh2:cf_role = "mesh_topology" ;
		Mesh2:topology_dimension = 2 ;
		Mesh2:long_name = "Topology data of 2D unstructured mesh" ;
		Mesh2:node_coordinates = "Mesh2_node_x Mesh2_node_y" ;
		Mesh2:edge_coordinates = "Mesh2_edge_x Mesh2_edge_y" ;
		Mesh2:face_coordinates = "Mesh2_face_x Mesh2_face_y" ;
		Mesh2:face_node_connectivity = "Mesh2_face_nodes" ;
		Mesh2:edge_node_connectivity = "Mesh2_edge_nodes" ;
		Mesh2:face_edge_connectivity = "Mesh2_face_edges" ;
		Mesh2:face_face_connectivity = "Mesh2_face_links" ;
		Mesh2:edge_face_connectivity = "Mesh2_edge_face_links" ;
	double Mesh2_node_x(nMesh2_node) ;
		Mesh2_node_x:units = "degrees_east" ;
		Mesh2_node_x:standard_name = "longitude" ;
		Mesh2_node_x:long_name = "Longitude of 2D mesh nodes." ;
	double Mesh2_node_y(nMesh2_node) ;
		Mesh2_node_y:units = "degrees_north" ;
		Mesh2_node_y:standard_name = "latitude" ;
		Mesh2_node_y:long_name = "Latitude of 2D mesh nodes." ;
	double Mesh2_edge_x(nMesh2_edge) ;
		Mesh2_edge_x:units = "degrees_east" ;
		Mesh2_edge_x:standard_name = "longitude" ;
		Mesh2_edge_x:long_name = "Characteristic longitude of 2D mesh edge (e.g. midpoint of the edge)." ;
	double Mesh2_edge_y(nMesh2_edge) ;
		Mesh2_edge_y:units = "degrees_north" ;
		Mesh2_edge_y:standard_name = "latitude" ;
		Mesh2_edge_y:long_name = "Characteristic latitude of 2D mesh edge (e.g. midpoint of the edge)." ;
	double Mesh2_face_x(nMesh2_face) ;
		Mesh2_face_x:units = "degrees_east" ;
		Mesh2_face_x:standard_name = "longitude" ;
		Mesh2_face_x:long_name = "Characteristics longitude of 2D mesh face." ;
	double Mesh2_face_y(nMesh2_face) ;
		Mesh2_face_y:units = "degrees_north" ;
		Mesh2_face_y:standard_name = "latitude" ;
		Mesh2_face_y:long_name = "Characteristics latitude of 2D mesh face." ;
	int Mesh2_face_nodes(nMesh2_face, Mesh2_face_N_nodes) ;
		Mesh2_face_nodes:long_name = "Maps every face to its corner nodes." ;
		Mesh2_face_nodes:cf_role = "face_node_connectivity" ;
		Mesh2_face_nodes:start_index = 1 ;
	int Mesh2_edge_nodes(nMesh2_edge, Mesh2_edge_N_nodes) ;
		Mesh2_edge_nodes:long_name = "Maps every edge to the two nodes that it connects." ;
		Mesh2_edge_nodes:cf_role = "edge_node_connectivity" ;
		Mesh2_edge_nodes:start_index = 1 ;
	int Mesh2_face_edges(nMesh2_face, Mesh2_face_N_edges) ;
		Mesh2_face_edges:long_name = "Maps every face to its edges." ;
		Mesh2_face_edges:cf_role = "face_edge_connectivity" ;
		Mesh2_face_edges:start_index = 1 ;
	int Mesh2_face_links(nMesh2_face, Mesh2_face_N_faces) ;
		Mesh2_face_links:long_name = "neighbor faces for faces" ;
		Mesh2_face_links:comment = "missing edges as well as missing neighbor faces are indicated using _FillValue" ;
		Mesh2_face_links:cf_role = "face_face_connectivity" ;
		Mesh2_face_links:start_index = 1 ;
	int Mesh2_edge_face_links(nMesh2_edge, Mesh2_edge_N_faces) ;
		Mesh2_edge_face_links:long_name = "neighbor faces for edges" ;
		Mesh2_edge_face_links:comment = "missing neighbor faces are indicated using _FillValue" ;
		Mesh2_edge_face_links:cf_role = "edge_face_connectivity" ;
		Mesh2_edge_face_links:start_index = 1 ;
	float datavar(Mesh2_layers, nMesh2_face) ;
		datavar:mesh = "Mesh2" ;
		datavar:location = "face" ;
		datavar:coordinates = "Mesh2_depth Mesh2_surface" ;
	double Mesh2_layers(Mesh2_layers) ;
		Mesh2_layers:axis = "Z" ;
		Mesh2_layers:units = "1" ;
		Mesh2_layers:standard_name = "ocean_sigma_coordinate" ;
		Mesh2_layers:long_name = "sigma at layer midpoints" ;
		Mesh2_layers:positive = "up" ;
		Mesh2_layers:formula_terms = "sigma: Mesh2_layers eta: Mesh2_surface depth: Mesh2_depth" ;
	double Mesh2_depth(nMesh2_face) ;
		Mesh2_depth:units = "m" ;
		Mesh2_depth:standard_name = "sea_floor_depth_below_geoid" ;
		Mesh2_depth:location = "face" ;
		Mesh2_depth:mesh = "Mesh2" ;
		Mesh2_depth:positive = "down" ;
	double Mesh2_surface(nMesh2_face) ;
		Mesh2_surface:units = "m" ;
		Mesh2_surface:standard_name = "sea_surface_height_above_geoid" ;
		Mesh2_surface:location = "face" ;
		Mesh2_surface:mesh = "Mesh2" ;
	double Mesh2_depth_0(nMesh2_face) ;
		Mesh2_depth_0:standard_name = "sea_floor_depth_below_geoid" ;
		Mesh2_depth_0:units = "m" ;
		Mesh2_depth_0:positive = "down" ;
		Mesh2_depth_0:mesh = "Mesh2" ;
		Mesh2_depth_0:location = "face" ;
	double Mesh2_surface_0(nMesh2_face) ;
		Mesh2_surface_0:standard_name = "sea_surface_height_above_geoid" ;
		Mesh2_surface_0:units = "m" ;
		Mesh2_surface_0:mesh = "Mesh2" ;
		Mesh2_surface_0:location = "face" ;

// global attributes:
		:Conventions = "CF-1.7" ;
}
