dimensions:
	bnds = 2 ;
	latitude = 73 ;
	pressure = 15 ;
variables:
	float geopotential_height(pressure, latitude) ;
		geopotential_height:_FillValue = 9.96921e+36f ;
		geopotential_height:standard_name = "geopotential_height" ;
		geopotential_height:units = "m" ;
		geopotential_height:um_stash_source = "m01s16i202" ;
		geopotential_height:cell_methods = "time: mean (interval: 4 hour)" ;
		geopotential_height:grid_mapping = "latitude_longitude" ;
		geopotential_height:coordinates = "forecast_period forecast_reference_time time" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	float pressure(pressure) ;
		pressure:axis = "Z" ;
		pressure:units = "hPa" ;
		pressure:long_name = "pressure" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	double forecast_period ;
		forecast_period:bounds = "forecast_period_bnds" ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	double forecast_period_bnds(bnds) ;
	double forecast_reference_time ;
		forecast_reference_time:units = "hours since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "360_day" ;
	double time ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(bnds) ;

// global attributes:
		:source = "Data from Met Office Unified Model" ;
		:Conventions = "CF-1.7" ;
}
