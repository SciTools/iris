dimensions:
	forecast_period = 4 ;
	latitude = 13 ;
	longitude = 10 ;
	bnds = 2 ;
variables:
	float unknown(forecast_period, latitude, longitude) ;
		unknown:cell_methods = "time: mean (interval: 1 hour)" ;
		unknown:grid_mapping = "latitude_longitude" ;
		unknown:coordinates = "forecast_reference_time height time" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:semi_major_axis = 6371229. ;
		latitude_longitude:semi_minor_axis = 6371229. ;
	int forecast_period(forecast_period) ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	double forecast_reference_time ;
		forecast_reference_time:units = "hours since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "360_day" ;
	double height ;
		height:units = "m" ;
		height:long_name = "height" ;
	double time(forecast_period) ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(forecast_period, bnds) ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:source = "Data from Met Office Unified Model" ;
}
