dimensions:
	time = UNLIMITED ; // (360 currently)
	bnds = 2 ;
	latitude = 73 ;
	longitude = 96 ;
variables:
	short air_temperature(time, latitude, longitude) ;
		air_temperature:scale_factor = 0.0024257504786326 ;
		air_temperature:add_offset = 261.648002426021 ;
		air_temperature:standard_name = "air_temperature" ;
		air_temperature:units = "K" ;
		air_temperature:um_stash_source = "m01s03i236" ;
		air_temperature:cell_methods = "time: maximum (interval: 1 hour)" ;
		air_temperature:grid_mapping = "latitude_longitude" ;
		air_temperature:coordinates = "forecast_period forecast_reference_time height" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	double forecast_period(time) ;
		forecast_period:bounds = "forecast_period_bnds" ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	double forecast_period_bnds(time, bnds) ;
	double forecast_reference_time ;
		forecast_reference_time:units = "hours since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "360_day" ;
	double height ;
		height:units = "m" ;
		height:standard_name = "height" ;
		height:positive = "up" ;
	float precipitation_flux(time, latitude, longitude) ;
		precipitation_flux:_FillValue = -1.e+30f ;
		precipitation_flux:standard_name = "precipitation_flux" ;
		precipitation_flux:units = "kg m-2 s-1" ;
		precipitation_flux:um_stash_source = "m01s05i216" ;
		precipitation_flux:cell_methods = "time: mean (interval: 1 hour)" ;
		precipitation_flux:grid_mapping = "latitude_longitude" ;
		precipitation_flux:coordinates = "forecast_period forecast_reference_time" ;
	ushort air_temperature_0(time, latitude, longitude) ;
		air_temperature_0:scale_factor = 0.0020141666756075 ;
		air_temperature_0:add_offset = 176.7872f ;
		air_temperature_0:standard_name = "air_temperature" ;
		air_temperature_0:units = "K" ;
		air_temperature_0:um_stash_source = "m01s03i236" ;
		air_temperature_0:cell_methods = "time: minimum (interval: 1 hour)" ;
		air_temperature_0:grid_mapping = "latitude_longitude" ;
		air_temperature_0:coordinates = "forecast_period forecast_reference_time height" ;

// global attributes:
		:source = "Data from Met Office Unified Model" ;
		:Conventions = "CF-1.5" ;
}
