dimensions:
	bnds = 2 ;
	site_number = 3 ;
	time = 240 ;
variables:
	float air_temperature(time, site_number) ;
		air_temperature:_FillValue = 9.96921e+36f ;
		air_temperature:standard_name = "air_temperature" ;
		air_temperature:units = "Celsius" ;
		air_temperature:um_stash_source = "m01s03i236" ;
		air_temperature:cell_methods = "time: mean" ;
		air_temperature:grid_mapping = "latitude_longitude" ;
		air_temperature:coordinates = "height latitude longitude" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	float time(time) ;
		time:axis = "T" ;
		time:units = "days since 0000-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	float site_number(site_number) ;
		site_number:units = "1" ;
		site_number:long_name = "site_number" ;
	double height ;
		height:units = "m" ;
		height:standard_name = "height" ;
	float latitude(site_number) ;
		latitude:bounds = "latitude_bnds" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	float latitude_bnds(site_number, bnds) ;
	float longitude(site_number) ;
		longitude:bounds = "longitude_bnds" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	float longitude_bnds(site_number, bnds) ;

// global attributes:
		:source = "Data from Met Office Unified Model" ;
		:Conventions = "CF-1.7" ;
}
