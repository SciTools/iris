dimensions:
	dim0 = 2 ;
	dim0_0 = 1 ;
	dim1 = 2 ;
	dim2 = 2 ;
variables:
	double temp(dim0, dim1) ;
		temp:standard_name = "surface_temperature" ;
		temp:units = "K" ;
		temp:history = "Team A won." ;
	double temp2(dim0_0, dim1, dim2) ;
		temp2:long_name = "Something Random" ;
		temp2:units = "K" ;
		temp2:history = "Team B won." ;

// global attributes:
		:Conventions = "CF-1.7" ;
}
