dimensions:
	latitude = 3 ;
	longitude = 4 ;
variables:
	int unknown(latitude, longitude) ;
		unknown:ukmo__process_flags = "X-derivative_(d/dx)" ;
		unknown:grid_mapping = "latitude_longitude" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	int latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	int longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;

// global attributes:
		:Conventions = "CF-1.7" ;
}
