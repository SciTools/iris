dimensions:
	bnds = 2 ;
	bnds_4 = 4 ;
	deptht = 31 ;
	dim2 = 148 ;
	dim3 = 180 ;
	time_counter = 1 ;
variables:
	float votemper(time_counter, deptht, dim2, dim3) ;
		votemper:standard_name = "sea_water_potential_temperature" ;
		votemper:long_name = "Temperature" ;
		votemper:units = "degC" ;
		votemper:cell_methods = "time_counter: mean" ;
		votemper:coordinates = "nav_lat nav_lon" ;
		votemper:cell_measures = "area: areat" ;
	float time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:units = "seconds since 0001-01-01 00:00:00" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "360_day" ;
		time_counter:time_origin = " 0001-JAN-01 00:00:00" ;
		time_counter:title = "Time" ;
	float deptht(deptht) ;
		deptht:axis = "Z" ;
		deptht:bounds = "deptht_bnds" ;
		deptht:units = "m" ;
		deptht:standard_name = "depth" ;
		deptht:long_name = "Vertical T levels" ;
		deptht:positive = "down" ;
		deptht:title = "deptht" ;
		deptht:valid_max = 5250.227f ;
		deptht:valid_min = 4.999938f ;
	double deptht_bnds(deptht, bnds) ;
	float nav_lat(dim2, dim3) ;
		nav_lat:bounds = "nav_lat_bnds" ;
		nav_lat:units = "degrees_north" ;
		nav_lat:standard_name = "latitude" ;
		nav_lat:long_name = "Latitude" ;
		nav_lat:nav_model = "Default grid" ;
		nav_lat:valid_max = 89.6139f ;
		nav_lat:valid_min = -78.19058f ;
	double nav_lat_bnds(dim2, dim3, bnds_4) ;
	float nav_lon(dim2, dim3) ;
		nav_lon:bounds = "nav_lon_bnds" ;
		nav_lon:units = "degrees_east" ;
		nav_lon:standard_name = "longitude" ;
		nav_lon:long_name = "Longitude" ;
		nav_lon:nav_model = "Default grid" ;
		nav_lon:valid_max = 180.f ;
		nav_lon:valid_min = -179.7507f ;
	double nav_lon_bnds(dim2, dim3, bnds_4) ;
	double areat(dim2, dim3) ;
		areat:units = "m2" ;
		areat:standard_name = "cell_area" ;
		areat:long_name = "area of grid cell" ;

// global attributes:
		:DOMAIN_DIM_N001 = "x" ;
		:DOMAIN_DIM_N002 = "y" ;
		:DOMAIN_DIM_N003 = "ncorners" ;
		:DOMAIN_DIM_N004 = "deptht" ;
		:DOMAIN_DIM_N005 = "ndepth_bounds" ;
		:DOMAIN_DIM_N006 = "time_counter" ;
		:DOMAIN_dimensions_ids = 1, 2 ;
		:DOMAIN_halo_size_end = 0, 0 ;
		:DOMAIN_halo_size_start = 0, 0 ;
		:DOMAIN_number = 0 ;
		:DOMAIN_number_total = 1 ;
		:DOMAIN_position_first = 1, 1 ;
		:DOMAIN_position_last = 182, 149 ;
		:DOMAIN_size_global = 182, 149 ;
		:DOMAIN_size_local = 182, 149 ;
		:DOMAIN_type = "box" ;
		:NCO = "4.0.8" ;
		:TimeStamp = "2008-SEP-09 11:18:37 GMT+0000" ;
		:file_name = "ORCA2_1d_00010101_00010101_grid_T_0000.nc" ;
		:history = "Mon Apr  2 10:25:46 2012: /project/ukmo/rhel6/nco/bin/ncks -v votemper,deptht_bounds,nav_lat,nav_lon,areat,latt_bounds,lont_bounds ORCA2_1d_00010101_00010101_grid_T_0000.nc votemper.nc" ;
		:interval_operation = 5760.f ;
		:interval_write = 86400.f ;
		:production = "An IPSL model" ;
		:short_name = "votemper" ;
		:Conventions = "CF-1.7" ;
}
