dimensions:
	bnds = 2 ;
	latitude = 3 ;
	longitude = 5 ;
	time = 4 ;
variables:
	byte climatology_test(time, latitude, longitude) ;
		climatology_test:long_name = "climatology test" ;
		climatology_test:units = "Kelvin" ;
		climatology_test:cell_methods = "time: mean over years" ;
	double time(time) ;
		time:axis = "T" ;
		time:climatology = "time_climatology" ;
		time:units = "days since 1970-01-01 00:00:00-00" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;
	double time_climatology(time, bnds) ;
	double latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "1" ;
		latitude:standard_name = "latitude" ;
	double longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "1" ;
		longitude:standard_name = "longitude" ;
}
