dimensions:
	bnds = 2 ;
	latitude = 73 ;
	longitude = 96 ;
	pressure = 15 ;
	time = 2 ;
variables:
	float geopotential_height(time, pressure, latitude, longitude) ;
		geopotential_height:standard_name = "geopotential_height" ;
		geopotential_height:units = "m" ;
		geopotential_height:um_stash_source = "m01s16i202" ;
		geopotential_height:cell_methods = "time: mean" ;
		geopotential_height:grid_mapping = "latitude_longitude" ;
		geopotential_height:coordinates = "forecast_period forecast_reference_time" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	float pressure(pressure) ;
		pressure:axis = "Z" ;
		pressure:units = "hPa" ;
		pressure:long_name = "pressure" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	double forecast_period(time) ;
		forecast_period:bounds = "forecast_period_bnds" ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	double forecast_period_bnds(time, bnds) ;
	double forecast_reference_time ;
		forecast_reference_time:units = "hours since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "360_day" ;

// global attributes:
		:source = "Data from Met Office Unified Model" ;
		:Conventions = "CF-1.5" ;
}
