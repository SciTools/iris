dimensions:
	dim0 = UNLIMITED ; // (1 currently)
	dim0_0 = UNLIMITED ; // (2 currently)
	dim1 = 2 ;
	dim2 = 2 ;
variables:
	double temp2(dim0, dim1, dim2) ;
		temp2:long_name = "Something Random" ;
		temp2:units = "K" ;
		temp2:fruit = "orange" ;
	double temp3(dim0_0, dim1, dim2) ;
		temp3:long_name = "Something Random" ;
		temp3:units = "K" ;
		temp3:fruit = "lemon" ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:foo = "bar" ;
		:fruit = "apple" ;
}
