dimensions:
	dim0 = 1 ;
variables:
	int64 unknown(dim0) ;

// global attributes:
		:Conventions = "CF-1.7" ;
}
