dimensions:
	bnds = 2 ;
variables:
	float air_potential_temperature ;
		air_potential_temperature:standard_name = "air_potential_temperature" ;
		air_potential_temperature:units = "K" ;
		air_potential_temperature:grid_mapping = "rotated_latitude_longitude" ;
		air_potential_temperature:coordinates = "forecast_period grid_latitude grid_longitude level_height model_level_number sigma surface_altitude time" ;
	int rotated_latitude_longitude ;
		rotated_latitude_longitude:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_latitude_longitude:longitude_of_prime_meridian = 0. ;
		rotated_latitude_longitude:earth_radius = 6371229. ;
		rotated_latitude_longitude:grid_north_pole_latitude = 37.5 ;
		rotated_latitude_longitude:grid_north_pole_longitude = 177.5 ;
		rotated_latitude_longitude:north_pole_grid_longitude = 0. ;
		rotated_latitude_longitude:crs_wkt = "GEOGCRS[\"unnamed\",BASEGEOGCRS[\"unknown\",DATUM[\"unknown\",ELLIPSOID[\"unknown\",6371229,0,LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]]],PRIMEM[\"Greenwich\",0,ANGLEUNIT[\"degree\",0.0174532925199433],ID[\"EPSG\",8901]]],DERIVINGCONVERSION[\"unknown\",METHOD[\"PROJ ob_tran o_proj=latlon\"],PARAMETER[\"o_lon_p\",0,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9122]]],PARAMETER[\"o_lat_p\",37.5,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9122]]],PARAMETER[\"lon_0\",357.5,ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9122]]]],CS[ellipsoidal,2],AXIS[\"longitude\",east,ORDER[1],ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9122]]],AXIS[\"latitude\",north,ORDER[2],ANGLEUNIT[\"degree\",0.0174532925199433,ID[\"EPSG\",9122]]]]" ;
	double forecast_period ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	float grid_latitude ;
		grid_latitude:bounds = "grid_latitude_bnds" ;
		grid_latitude:units = "degrees" ;
		grid_latitude:standard_name = "grid_latitude" ;
	float grid_latitude_bnds(bnds) ;
	float grid_longitude ;
		grid_longitude:bounds = "grid_longitude_bnds" ;
		grid_longitude:units = "degrees" ;
		grid_longitude:standard_name = "grid_longitude" ;
	float grid_longitude_bnds(bnds) ;
	float level_height ;
		level_height:bounds = "level_height_bnds" ;
		level_height:units = "m" ;
		level_height:long_name = "level_height" ;
		level_height:positive = "up" ;
		level_height:standard_name = "atmosphere_hybrid_height_coordinate" ;
		level_height:axis = "Z" ;
		level_height:formula_terms = "a: level_height b: sigma orog: surface_altitude" ;
	float level_height_bnds(bnds) ;
	int model_level_number ;
		model_level_number:units = "1" ;
		model_level_number:standard_name = "model_level_number" ;
		model_level_number:positive = "up" ;
	float sigma ;
		sigma:bounds = "sigma_bnds" ;
		sigma:units = "1" ;
		sigma:long_name = "sigma" ;
	float sigma_bnds(bnds) ;
	float surface_altitude ;
		surface_altitude:units = "m" ;
		surface_altitude:standard_name = "surface_altitude" ;
	double time ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;

// global attributes:
		:source = "Iris test case" ;
		:Conventions = "CF-1.7" ;
}
