dimensions:
	bnds = 2 ;
	latitude = 3 ;
	longitude = 5 ;
	time = 4 ;
variables:
	byte climatology_test(time, latitude, longitude) ;
		climatology_test:long_name = "climatology test" ;
		climatology_test:units = "Kelvin" ;
		climatology_test:cell_methods = "time: mean over years" ;
	double time(time) ;
		time:axis = "T" ;
		time:units = "days since 1970-01-01 00:00:00-00" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;
		time:climatology = "time_climatology" ;
	double latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "1" ;
		latitude:standard_name = "latitude" ;
	double longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "1" ;
		longitude:standard_name = "longitude" ;
	double time_climatology(time, bnds) ;

// global attributes:
		:Conventions = "CF-1.5" ;
data:

 climatology_test =
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0 ;

 time = 11332, 11333, 11334, 11335 ;

 latitude = 0, 30, 60 ;

 longitude = -25, -12.5, 0, 12.5, 25 ;

 time_climatology =
  11332, 14984,
  11333, 14985,
  11334, 14986,
  11335, 14987 ;
}
