dimensions:
	dim0 = 4 ;
	dim1 = 5 ;
	string6 = 6 ;
variables:
	double unknown(dim0, dim1) ;
		unknown:coordinates = "unknown_scalar" ;
	double dim0(dim0) ;
		dim0:units = "1" ;
	double dim1(dim1) ;
		dim1:units = "m" ;
	char unknown_scalar(string6) ;

// global attributes:
		:Conventions = "CF-1.7" ;
}
