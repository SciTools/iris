dimensions:
	bnds = 2 ;
	depth = 20 ;
	grid_latitude = 143 ;
	pseudo_level = 4 ;
	time = 4 ;
variables:
	float unknown(pseudo_level, time, depth, grid_latitude) ;
		unknown:_FillValue = 9.96921e+36f ;
		unknown:um_stash_source = "m02s00i???" ;
		unknown:cell_methods = "time: mean" ;
		unknown:grid_mapping = "rotated_latitude_longitude" ;
		unknown:coordinates = "forecast_period forecast_reference_time" ;
	int rotated_latitude_longitude ;
		rotated_latitude_longitude:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_latitude_longitude:longitude_of_prime_meridian = 0. ;
		rotated_latitude_longitude:earth_radius = 6371229. ;
		rotated_latitude_longitude:grid_north_pole_latitude = 0. ;
		rotated_latitude_longitude:grid_north_pole_longitude = 0. ;
		rotated_latitude_longitude:north_pole_grid_longitude = 0. ;
	int pseudo_level(pseudo_level) ;
		pseudo_level:units = "1" ;
		pseudo_level:long_name = "pseudo_level" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	float depth(depth) ;
		depth:axis = "Z" ;
		depth:units = "m" ;
		depth:standard_name = "depth" ;
		depth:positive = "down" ;
	float grid_latitude(grid_latitude) ;
		grid_latitude:axis = "Y" ;
		grid_latitude:units = "degrees" ;
		grid_latitude:standard_name = "grid_latitude" ;
	double forecast_period(time) ;
		forecast_period:bounds = "forecast_period_bnds" ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	double forecast_period_bnds(time, bnds) ;
	double forecast_reference_time ;
		forecast_reference_time:units = "hours since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "360_day" ;

// global attributes:
		:source = "Data from Met Office Unified Model" ;
		:Conventions = "CF-1.5" ;
}
