dimensions:
	depth = UNLIMITED ; // (20 currently)
	time = 16 ;
variables:
	float unknown(depth, time) ;
		unknown:_FillValue = 9.96921e+36f ;
		unknown:um_stash_source = "m??s44i101" ;
		unknown:cell_methods = "time: mean (interval: 24 hour)" ;
	float depth(depth) ;
		depth:axis = "Z" ;
		depth:units = "m" ;
		depth:standard_name = "depth" ;
		depth:positive = "down" ;
	float time(time) ;
		time:axis = "T" ;
		time:units = "days since 0000-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;

// global attributes:
		:source = "Data from Met Office Unified Model" ;
		:Conventions = "CF-1.5" ;
}
