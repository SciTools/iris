dimensions:
	depth = UNLIMITED ; // (20 currently)
	bnds = 2 ;
	latitude = 73 ;
variables:
	float unknown(depth, latitude) ;
		unknown:_FillValue = -1.e+30f ;
		unknown:ukmo__um_stash_source = "m??s44i101" ;
		unknown:ukmo__process_flags = "Mean_over_an_ensemble_of_parallel_runs Time_mean_field" ;
		unknown:grid_mapping = "latitude_longitude" ;
		unknown:coordinates = "forecast_period forecast_reference_time time" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:semi_major_axis = 6371229. ;
		latitude_longitude:semi_minor_axis = 6371229. ;
	float depth(depth) ;
		depth:axis = "Z" ;
		depth:units = "m" ;
		depth:standard_name = "depth" ;
		depth:positive = "down" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	int forecast_period ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	double forecast_reference_time ;
		forecast_reference_time:units = "hours since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "360_day" ;
	double time ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(bnds) ;

// global attributes:
		:source = "Data from Met Office Unified Model" ;
		:Conventions = "CF-1.5" ;
}
