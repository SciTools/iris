dimensions:
	pseudo_level = UNLIMITED ; // (4 currently)
	bnds = 2 ;
	latitude = 143 ;
	longitude = 1 ;
	time = 4 ;
variables:
	float northward_ocean_heat_transport(pseudo_level, time, latitude, longitude) ;
		northward_ocean_heat_transport:_FillValue = -1.e+30f ;
		northward_ocean_heat_transport:standard_name = "northward_ocean_heat_transport" ;
		northward_ocean_heat_transport:units = "PW" ;
		northward_ocean_heat_transport:ukmo__um_stash_source = "m02s30i211" ;
		northward_ocean_heat_transport:source = "Data from Met Office Unified Model" ;
		northward_ocean_heat_transport:cell_methods = "time: mean" ;
		northward_ocean_heat_transport:grid_mapping = "latitude_longitude" ;
		northward_ocean_heat_transport:coordinates = "forecast_period forecast_reference_time" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:semi_major_axis = 6371229. ;
		latitude_longitude:semi_minor_axis = 6371229. ;
	int pseudo_level(pseudo_level) ;
		pseudo_level:units = "1" ;
		pseudo_level:long_name = "pseudo_level" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	int forecast_period(time) ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	double forecast_reference_time ;
		forecast_reference_time:units = "hours since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "360_day" ;

// global attributes:
		:Conventions = "CF-1.5" ;
}
