dimensions:
	bnds = 2 ;
	grid_latitude = 100 ;
	grid_longitude = 100 ;
	model_level_number = 70 ;
	time = 6 ;
variables:
	float air_potential_temperature(time, model_level_number, grid_latitude, grid_longitude) ;
		air_potential_temperature:standard_name = "air_potential_temperature" ;
		air_potential_temperature:units = "K" ;
		air_potential_temperature:grid_mapping = "rotated_latitude_longitude" ;
		air_potential_temperature:coordinates = "forecast_period level_height level_pressure sigma surface_air_pressure surface_altitude unknown_scalar" ;
	int rotated_latitude_longitude ;
		rotated_latitude_longitude:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_latitude_longitude:longitude_of_prime_meridian = 0. ;
		rotated_latitude_longitude:earth_radius = 6371229. ;
		rotated_latitude_longitude:grid_north_pole_latitude = 37.5 ;
		rotated_latitude_longitude:grid_north_pole_longitude = 177.5 ;
		rotated_latitude_longitude:north_pole_grid_longitude = 0. ;
	double time(time) ;
		time:axis = "T" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;
	int model_level_number(model_level_number) ;
		model_level_number:axis = "Z" ;
		model_level_number:units = "1" ;
		model_level_number:standard_name = "model_level_number" ;
		model_level_number:positive = "up" ;
	float grid_latitude(grid_latitude) ;
		grid_latitude:axis = "Y" ;
		grid_latitude:bounds = "grid_latitude_bnds" ;
		grid_latitude:units = "degrees" ;
		grid_latitude:standard_name = "grid_latitude" ;
	float grid_latitude_bnds(grid_latitude, bnds) ;
	float grid_longitude(grid_longitude) ;
		grid_longitude:axis = "X" ;
		grid_longitude:bounds = "grid_longitude_bnds" ;
		grid_longitude:units = "degrees" ;
		grid_longitude:standard_name = "grid_longitude" ;
	float grid_longitude_bnds(grid_longitude, bnds) ;
	double forecast_period ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	float level_height(model_level_number) ;
		level_height:bounds = "level_height_bnds" ;
		level_height:units = "m" ;
		level_height:long_name = "level_height" ;
		level_height:positive = "up" ;
		level_height:standard_name = "atmosphere_hybrid_height_coordinate" ;
		level_height:axis = "Z" ;
		level_height:formula_terms = "a: level_height b: sigma orog: surface_altitude" ;
	float level_height_bnds(model_level_number, bnds) ;
	double level_pressure ;
		level_pressure:units = "hPa" ;
		level_pressure:long_name = "level_pressure" ;
		level_pressure:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate" ;
		level_pressure:axis = "Z" ;
		level_pressure:formula_terms = "ap: level_pressure b: unknown_scalar ps: surface_air_pressure" ;
	double unknown_scalar ;
		unknown_scalar:units = "1" ;
		unknown_scalar:long_name = "other sigma" ;
	float sigma(model_level_number) ;
		sigma:bounds = "sigma_bnds" ;
		sigma:units = "1" ;
		sigma:long_name = "sigma" ;
	float sigma_bnds(model_level_number, bnds) ;
	double surface_air_pressure ;
		surface_air_pressure:units = "hPa" ;
		surface_air_pressure:long_name = "surface_air_pressure" ;
	float surface_altitude(grid_latitude, grid_longitude) ;
		surface_altitude:units = "m" ;
		surface_altitude:standard_name = "surface_altitude" ;

// global attributes:
		:source = "Iris test case" ;
		:Conventions = "CF-1.5" ;
}
