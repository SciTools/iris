dimensions:
	dim0 = UNLIMITED ; // (2 currently)
	dim0_0 = UNLIMITED ; // (1 currently)
	dim1 = 2 ;
	dim2 = 2 ;
variables:
	double temp(dim0, dim1) ;
		temp:standard_name = "surface_temperature" ;
		temp:units = "K" ;
		temp:foo = "bar" ;
	double temp2(dim0_0, dim1, dim2) ;
		temp2:long_name = "Something Random" ;
		temp2:units = "K" ;
		temp2:foo = "orange" ;

// global attributes:
		:Conventions = "CF-1.5" ;
}
