dimensions:
	grid_latitude = 2 ;
	grid_longitude = 2 ;
	latitude = 2 ;
	latitude_0 = 2 ;
	longitude = 2 ;
	longitude_0 = 2 ;
variables:
	int64 air_temperature(longitude, latitude) ;
		air_temperature:standard_name = "air_temperature" ;
		air_temperature:grid_mapping = "latitude_longitude" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	int64 longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "1" ;
	int64 latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "1" ;
	int64 air_temperature_0(longitude_0, latitude_0) ;
		air_temperature_0:standard_name = "air_temperature" ;
		air_temperature_0:grid_mapping = "latitude_longitude_0" ;
	int latitude_longitude_0 ;
		latitude_longitude_0:grid_mapping_name = "latitude_longitude_0" ;
		latitude_longitude_0:longitude_of_prime_meridian = 0. ;
		latitude_longitude_0:earth_radius = 6371228. ;
	int64 longitude_0(longitude_0) ;
		longitude_0:axis = "X" ;
		longitude_0:units = "degrees_east" ;
		longitude_0:standard_name = "longitude" ;
		longitude_0:long_name = "2" ;
	int64 latitude_0(latitude_0) ;
		latitude_0:axis = "Y" ;
		latitude_0:units = "degrees_north" ;
		latitude_0:standard_name = "latitude" ;
		latitude_0:long_name = "2" ;
	int64 air_temperature_1(grid_longitude, grid_latitude) ;
		air_temperature_1:standard_name = "air_temperature" ;
		air_temperature_1:grid_mapping = "rotated_latitude_longitude" ;
	int rotated_latitude_longitude ;
		rotated_latitude_longitude:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_latitude_longitude:grid_north_pole_latitude = 30. ;
		rotated_latitude_longitude:grid_north_pole_longitude = 30. ;
		rotated_latitude_longitude:north_pole_grid_longitude = 0. ;
	int64 grid_longitude(grid_longitude) ;
		grid_longitude:axis = "X" ;
		grid_longitude:units = "degrees" ;
		grid_longitude:standard_name = "grid_longitude" ;
		grid_longitude:long_name = "3" ;
	int64 grid_latitude(grid_latitude) ;
		grid_latitude:axis = "Y" ;
		grid_latitude:units = "degrees" ;
		grid_latitude:standard_name = "grid_latitude" ;
		grid_latitude:long_name = "3" ;

// global attributes:
		:Conventions = "CF-1.7" ;
}
