dimensions:
	bnds = 2 ;
	dim0 = 3 ;
	dim1 = 4 ;
variables:
	float air_pressure_anomaly(dim0, dim1) ;
		air_pressure_anomaly:standard_name = "air_pressure_anomaly" ;
	float dim0(dim0) ;
		dim0:bounds = "dim0_bnds" ;
		dim0:units = "1" ;
	float dim0_bnds(dim0, bnds) ;
}
