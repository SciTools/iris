dimensions:
	grid_latitude = 9 ;
	grid_longitude = 11 ;
	time = 7 ;
variables:
	int64 air_potential_temperature(time, grid_latitude, grid_longitude) ;
		air_potential_temperature:standard_name = "air_potential_temperature" ;
		air_potential_temperature:units = "K" ;
		air_potential_temperature:grid_mapping = "rotated_latitude_longitude" ;
		air_potential_temperature:coordinates = "air_pressure forecast_period" ;
		air_potential_temperature:ancillary_variables = "latlon_refs" ;
	int rotated_latitude_longitude ;
		rotated_latitude_longitude:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_latitude_longitude:longitude_of_prime_meridian = 0. ;
		rotated_latitude_longitude:earth_radius = 6371229. ;
		rotated_latitude_longitude:grid_north_pole_latitude = 37.5 ;
		rotated_latitude_longitude:grid_north_pole_longitude = 177.5 ;
		rotated_latitude_longitude:north_pole_grid_longitude = 0. ;
	double time(time) ;
		time:axis = "T" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;
	double grid_latitude(grid_latitude) ;
		grid_latitude:axis = "Y" ;
		grid_latitude:units = "degrees" ;
		grid_latitude:standard_name = "grid_latitude" ;
	double grid_longitude(grid_longitude) ;
		grid_longitude:axis = "X" ;
		grid_longitude:units = "degrees" ;
		grid_longitude:standard_name = "grid_longitude" ;
	double air_pressure ;
		air_pressure:units = "Pa" ;
		air_pressure:standard_name = "air_pressure" ;
	double forecast_period(time) ;
		forecast_period:units = "hours" ;
		forecast_period:standard_name = "forecast_period" ;
	double latlon_refs(grid_latitude, grid_longitude) ;
		latlon_refs:units = "s" ;
		latlon_refs:long_name = "latlon_refs" ;
	int64 alternate_data(time, grid_latitude, grid_longitude) ;
		alternate_data:long_name = "alternate_data" ;
		alternate_data:units = "m" ;
		alternate_data:grid_mapping = "rotated_latitude_longitude" ;
		alternate_data:coordinates = "air_pressure forecast_period" ;
		alternate_data:ancillary_variables = "latlon_refs_0" ;
	double latlon_refs_0(grid_latitude, grid_longitude) ;
		latlon_refs_0:units = "s" ;
		latlon_refs_0:long_name = "latlon_refs" ;

// global attributes:
		:source = "Iris test case" ;
		:Conventions = "CF-1.7" ;
}
